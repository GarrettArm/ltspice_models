PENTODE CHARACTERISTIC CURVES

* SET THESE TWO PARAMETERS FOR MODE (PENTODE, UL, TRIODE)
.PARAM TRIMODE = 40      ; % TRIODE MODE (0=PENTODE; 40=UL; 100=TRI...)
.PARAM VG2NOM = 450      ; NOMINAL VALUE OF GRID 2 VOLTAGE.
.STEP LIN VG1 0 -75 -10 ; 15 -75 -15  ; STEPS FOR PLATE CURVES

.PARAM T1 = {TRIMODE/100}, T2 = {1-T1}  ; FRACTION TRIODE MODE...
V_P 101 0 400  ; PLATE VOLTAGE
VP 101 1 0     ; DUMMY V SOURCE FOR POSITIVE PLATE CURRENT PLOT.
EG2 102 0 VALUE={VG2NOM*T2+T1*V(101,0)}  ; GRID 2 VOLTAGE 
VG2 102 4 0    ; FOR G2 CURRENT MEAS.
VG1 2 0 0      ; CONTROL GRID VOLTAGE
VC  3 0 0    ; FOR CATHODE CURRENT MEAS.
X1 1 2 3 4 6550  ; P G1 C G2
.DC LIN V_P  0 600 5    ; VB IS THE SUPPLY VOLTAGE.  I(VB) IS OUTPUT.
.PROBE I(VC) I(VP) I(VG2) I(VG1)
.OPTIONS NOPAGE LIBRARY
.LIB C:\PSPICE\WORK\TUBE.LIB
.END 